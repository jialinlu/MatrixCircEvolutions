*g_0_i_2_subckt.cir 
.SUBCKT HOT_CIRCUIT 5 28 3 vsupp vsupn 
R_0 1 2 94569.7042149 
R_2 3 4 6251290.57634 
x_4 5 5 7 par3pnp 
x_7 5 5 2 par3pnp 
q_10 11 5 11 BC308B 
xmn_13 3 3 11 0 submodn w=1.57962582294e-06 l=3.1106741486e-06 m=1 
xmn_16 17 4 1 0 submodn w=6.60809345571e-06 l=4.01068321349e-07 m=1 
xmn_19 3 3 3 0 submodn w=2.37462376849e-05 l=1.85723725489e-06 m=1 
xmn_22 23 3 17 0 submodn w=9.46481964864e-05 l=3.99349312183e-06 m=1 
xmp_25 26 27 28 vdd submodp w=2.1574867072e-06 l=2.72520969647e-06 m=1 
xmp_28 27 27 28 vdd submodp w=4.13143976161e-05 l=1.49836419629e-06 m=1 
xmp_31 3 23 26 vdd submodp w=7.09373980507e-05 l=1.16566221989e-06 m=1 
xmp_34 23 23 27 vdd submodp w=8.86444458606e-05 l=2.01256520897e-07 m=1 
xmp_37 38 27 28 vdd submodp w=5.18765948507e-05 l=4.35566959303e-07 m=1 
xmp_40 3 23 38 vdd submodp w=9.67772538715e-05 l=3.58796700611e-06 m=1 

*Convergence-aid resistors:
R_40 1 0 1e9 
R_41 2 0 1e9 
R_42 3 0 1e9 
R_43 4 0 1e9 
R_44 5 0 1e9 
R_77 38 0 1e9 
R_46 7 0 1e9 
R_50 11 0 1e9 
R_56 17 0 1e9 
R_62 23 0 1e9 
R_65 26 0 1e9 
R_66 27 0 1e9 
R_67 28 0 1e9 
.ends
