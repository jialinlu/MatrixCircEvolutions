*g_0_i_3_subckt.cir 
.SUBCKT HOT_CIRCUIT 2 28 3 vsupp vsupn 
R_0 1 2 146919.643966 
*R_2 3 3 12028.2057683 
*x_4 2 2 2 par3pnp 
*x_7 2 2 2 par3pnp 
*q_10 2 2 2 BC308B 
xmn_13 14 14 2 0 submodn w=4.09245405702e-07 l=3.93456807092e-07 m=1 
xmn_16 17 3 1 0 submodn w=3.91358723909e-06 l=3.51065677843e-07 m=1 
xmn_19 3 3 14 0 submodn w=3.37766190787e-06 l=3.73004775634e-06 m=1 
xmn_22 23 3 17 0 submodn w=7.2082766889e-05 l=1.51249302224e-06 m=1 
xmp_25 26 27 28 vdd submodp w=8.07305386921e-05 l=3.98587004416e-06 m=1 
xmp_28 27 27 28 vdd submodp w=7.27062166717e-05 l=1.49510190623e-06 m=1 
xmp_31 3 23 26 vdd submodp w=7.91673584347e-05 l=1.57089827297e-06 m=1 
xmp_34 23 23 27 vdd submodp w=8.79523882625e-05 l=2.07252963529e-07 m=1 
xmp_37 38 27 28 vdd submodp w=3.44058583244e-05 l=3.12182400562e-06 m=1 
xmp_40 3 23 38 vdd submodp w=4.84344911818e-05 l=3.74885457199e-06 m=1 

*Convergence-aid resistors:
R_40 1 0 1e9 
R_41 2 0 1e9 
R_42 3 0 1e9 
R_77 38 0 1e9 
R_53 14 0 1e9 
R_56 17 0 1e9 
R_62 23 0 1e9 
R_65 26 0 1e9 
R_66 27 0 1e9 
R_67 28 0 1e9 
.ends
