*g_0_i_0_subckt.cir 
.SUBCKT HOT_CIRCUIT 5 22 3 vsupp vsupn 
R_0 1 2 94569.7042149 
R_2 3 4 9446841.84997 
x_4 5 5 7 par3pnp 
x_7 5 5 2 par3pnp 
q_10 11 5 11 BC308B 
xmn_13 3 3 11 0 submodn w=1.57962582294e-06 l=2.97908882518e-06 m=1 
xmn_16 17 4 1 0 submodn w=1.36929320905e-05 l=4.59265712853e-07 m=1 
xmn_19 3 3 22 0 submodn w=7.07715100993e-05 l=3.29807718758e-06 m=1 
xmn_22 23 3 17 0 submodn w=9.65918952381e-05 l=1.31427848365e-06 m=1 
xmp_25 26 27 22 vdd submodp w=2.1574867072e-06 l=3.82372578463e-06 m=1 
xmp_28 27 27 22 vdd submodp w=4.02921173217e-05 l=1.49836419629e-06 m=1 
xmp_31 3 23 26 vdd submodp w=8.94767601645e-05 l=2.83696171269e-06 m=1 
xmp_34 23 23 27 vdd submodp w=5.73118515408e-05 l=2.01256520897e-07 m=1 
xmp_37 38 27 22 vdd submodp w=5.1152962751e-05 l=4.35566959303e-07 m=1 
xmp_40 3 23 38 vdd submodp w=9.56884969812e-05 l=3.83904970969e-06 m=1 

*Convergence-aid resistors:
R_40 1 0 1e9 
R_41 2 0 1e9 
R_42 3 0 1e9 
R_43 4 0 1e9 
R_44 5 0 1e9 
R_77 38 0 1e9 
R_46 7 0 1e9 
R_50 11 0 1e9 
R_56 17 0 1e9 
R_61 22 0 1e9 
R_62 23 0 1e9 
R_65 26 0 1e9 
R_66 27 0 1e9 
.ends
