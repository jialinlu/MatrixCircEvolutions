*g_0_i_0_subckt.cir 
.SUBCKT HOT_CIRCUIT 6 3 1 vsupp vsupn 
*R_0 1 1 2027122.49721 
*R_2 3 3 6915196.70387 
x_4 5 6 7 par3pnp 
x_7 3 3 1 par3pnp 
q_10 1 7 1 BC308B 
xmn_13 14 14 3 0 submodn w=4.89914957729e-05 l=1.34130937112e-06 m=1 
xmn_16 17 14 19 0 submodn w=2.43995028895e-05 l=1.54241640107e-06 m=1 
xmn_19 6 17 22 0 submodn w=5.18774591163e-05 l=3.34748685773e-06 m=1 
xmn_22 3 19 22 0 submodn w=8.87423896636e-05 l=3.13662297439e-06 m=1 
xmp_25 19 3 3 vdd submodp w=8.98254857034e-05 l=1.5550195994e-06 m=1 
xmp_28 14 5 14 vdd submodp w=2.67161210949e-05 l=2.80233506941e-06 m=1 
xmp_31 22 33 1 vdd submodp w=3.70637756516e-05 l=1.78189001685e-06 m=1 
xmp_34 14 22 14 vdd submodp w=6.62393791721e-05 l=1.23328551128e-06 m=1 
xmp_37 3 6 22 vdd submodp w=2.03996171556e-06 l=3.25813363966e-06 m=1 
xmp_40 7 3 3 vdd submodp w=3.60204833558e-05 l=2.57851056581e-06 m=1 

*Convergence-aid resistors:
R_35 1 0 1e9 
R_37 3 0 1e9 
R_39 5 0 1e9 
R_40 6 0 1e9 
R_41 7 0 1e9 
R_48 14 0 1e9 
R_51 17 0 1e9 
R_53 19 0 1e9 
R_56 22 0 1e9 
R_67 33 0 1e9 
.ends
