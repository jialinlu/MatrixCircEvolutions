*g_0_i_0_subckt.cir 
.SUBCKT HOT_CIRCUIT 2 22 14 vsupp vsupn 
R_0 1 2 69537.3985911 
R_2 3 4 30460.859214 
x_4 2 6 6 par3pnp 
x_7 2 3 6 par3pnp 
q_10 2 2 13 BC308B 
xmn_13 14 14 13 0 submodn w=1.80081798521e-07 l=2.23044678459e-06 m=1 
xmn_16 17 14 1 0 submodn w=1.33474214669e-05 l=3.39035075657e-07 m=1 
xmn_19 14 14 22 0 submodn w=9.07000614905e-05 l=3.47329692752e-06 m=1 
xmn_22 23 14 17 0 submodn w=9.99999970806e-05 l=1.19096216018e-06 m=1 
xmp_25 26 27 22 vdd submodp w=9.99999999812e-05 l=7.17033299916e-07 m=1 
xmp_28 27 27 22 vdd submodp w=2.61490239874e-05 l=2.17968621926e-07 m=1 
xmp_31 14 23 26 vdd submodp w=5.80652529759e-05 l=3.99999870618e-06 m=1 
xmp_34 23 23 27 vdd submodp w=6.65959000577e-05 l=1.98758423858e-07 m=1 
xmp_37 1 14 1 vdd submodp w=9.97480124893e-05 l=3.42866361039e-06 m=1 
xmp_40 1 6 6 vdd submodp w=9.99988657149e-05 l=2.01131245279e-07 m=1 

*Convergence-aid resistors:
R_29 1 0 1e9 
R_30 2 0 1e9 
R_31 3 0 1e9 
R_32 4 0 1e9 
R_34 6 0 1e9 
R_41 13 0 1e9 
R_42 14 0 1e9 
R_45 17 0 1e9 
R_50 22 0 1e9 
R_51 23 0 1e9 
R_54 26 0 1e9 
R_55 27 0 1e9 
.ends
