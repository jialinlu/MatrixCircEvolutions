*g_0_i_0_subckt.cir 
.SUBCKT HOT_CIRCUIT 2 28 3 vsupp vsupn 
R_0 1 2 207900.825134 
*R_2 3 3 6591792.58601 
x_4 2 2 7 par3pnp 
*x_7 2 2 2 par3pnp 
*q_10 2 2 2 BC308B 
xmn_13 14 14 2 0 submodn w=5.04388340215e-07 l=2.09367463788e-06 m=1 
xmn_16 17 3 1 0 submodn w=4.40540899757e-06 l=6.42222954358e-07 m=1 
xmn_19 3 3 14 0 submodn w=2.00589376677e-06 l=3.08874280763e-06 m=1 
xmn_22 23 3 17 0 submodn w=9.76540531057e-05 l=2.51590886506e-06 m=1 
xmp_25 26 27 28 vdd submodp w=9.62539781304e-05 l=8.38526952395e-07 m=1 
xmp_28 27 27 28 vdd submodp w=2.48187580347e-05 l=2.4696889193e-07 m=1 
xmp_31 3 23 26 vdd submodp w=9.9676582845e-05 l=3.91933708008e-06 m=1 
xmp_34 23 23 27 vdd submodp w=6.33831262965e-05 l=1.92704750062e-07 m=1 
xmp_37 38 27 28 vdd submodp w=8.53179022675e-05 l=3.66747650114e-06 m=1 
xmp_40 3 23 38 vdd submodp w=6.03206589488e-05 l=3.99669547282e-06 m=1 

*Convergence-aid resistors:
R_40 1 0 1e9 
R_41 2 0 1e9 
R_42 3 0 1e9 
R_77 38 0 1e9 
R_46 7 0 1e9 
R_53 14 0 1e9 
R_56 17 0 1e9 
R_62 23 0 1e9 
R_65 26 0 1e9 
R_66 27 0 1e9 
R_67 28 0 1e9 
.ends
