*g_1234_i_1234_subckt.cir 
.SUBCKT HOT_CIRCUIT 2 28 3 vsupp vsupn 
R_0 1 2 94569.7042149 
*R_2 3 3 4786003.90052 
x_4 2 2 7 par3pnp 
*x_7 2 2 2 par3pnp 
*q_10 2 2 2 BC308B 
xmn_13 14 14 2 0 submodn w=2.69531420894e-07 l=2.84493828712e-06 m=1 
xmn_16 17 3 1 0 submodn w=5.62643196646e-06 l=2.5972722024e-07 m=1 
xmn_19 3 3 14 0 submodn w=2.39522191933e-05 l=2.49464572401e-07 m=1 
xmn_22 23 3 17 0 submodn w=9.47189144413e-05 l=3.20236118445e-07 m=1 
xmp_25 2 2 28 vdd submodp w=2.1574867072e-06 l=3.66745611268e-06 m=1 
xmp_28 23 23 28 vdd submodp w=5.17762084718e-05 l=1.76854752919e-06 m=1 
xmp_31 3 23 34 vdd submodp w=9.93382504472e-05 l=1.89657483446e-07 m=1 
xmp_34 23 23 23 vdd submodp w=2.80190311935e-05 l=5.27569340482e-07 m=1 
xmp_37 34 23 28 vdd submodp w=3.46744021546e-05 l=3.99923671553e-06 m=1 
xmp_40 41 23 34 vdd submodp w=3.58780531207e-05 l=2.47721426019e-06 m=1 

*Convergence-aid resistors:
R_43 1 0 1e9 
R_44 2 0 1e9 
R_45 3 0 1e9 
R_49 7 0 1e9 
R_83 41 0 1e9 
R_76 34 0 1e9 
R_56 14 0 1e9 
R_59 17 0 1e9 
R_65 23 0 1e9 
R_70 28 0 1e9 
.ends
